package timing_parameters;
 
parameter tRC      = 115;
parameter tRAS      = 76;
parameter tRRD_L      = 12;
parameter tRRD_S      = 8;
parameter tRP      = 39;
parameter tRFC      = 295; // 295ns
parameter tCWD        = 38;
parameter tCAS        = 40;
parameter tRCD      = 39;
parameter tWR      = 30;
parameter tRTP      = 18;
parameter tCCD_L      = 12;
parameter tCCD_S      = 8;
parameter tCCD_L_WR   = 48;
parameter tCCD_S_WR   = 8;
parameter tBURST      = 8;
parameter tCCD_L_RTW  = 16;
parameter tCCD_S_RTW  = 16;
parameter tCCD_L_WTR  = 70;
parameter tCCD_S_WTR  = 52;
 

endpackage
