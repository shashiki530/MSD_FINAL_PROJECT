//////////////////
controller
