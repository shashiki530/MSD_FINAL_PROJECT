package timing_parameters;
 
parameter tRC 	      = 2*115;
parameter tRAS 	      = 2* 76; 
parameter tRRD_L      = 2* 12; 
parameter tRRD_S      = 2* 8; 
parameter tRP 	      = 2* 39; 
parameter tRFC 	      = 2* 295; // 295ns 
parameter tCWL        = 2* 38; 
parameter tCAS        = 2* 40; 
parameter tRCD 	      = 2* 39; 
parameter tWR 	      = 2* 30; 
parameter tRTP 	      = 2* 18; 
parameter tCCD_L      = 2* 12; 
parameter tCCD_S      = 2* 8; 
parameter tCCD_L_WR   = 2* 48; 
parameter tCCD_S_WR   = 2* 8; 
parameter tBURST      = 2* 8; 
parameter tCCD_L_RTW  = 2* 16; 
parameter tCCD_S_RTW  = 2* 16; 
parameter tCCD_L_WTR  = 2* 70; 
parameter tCCD_S_WTR  = 2* 52; 
 

endpackage

